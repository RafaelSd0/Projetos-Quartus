library verilog;
use verilog.vl_types.all;
entity Teste_vlg_vec_tst is
end Teste_vlg_vec_tst;
