library verilog;
use verilog.vl_types.all;
entity Teste_vlg_check_tst is
    port(
        o               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Teste_vlg_check_tst;
